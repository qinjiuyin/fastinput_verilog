module fastinput (
    input rst,
    input clk,

    output tx,
    input rx
);

endmodule
